module fsm_b (state, odd , even, terminal, pause, restart, clk, rst, goto_third, Out1, Out2);
	
	input pause, restart, clk, rst, goto_third;
	output reg [2:0] Out1, Out2;
	output odd, even, terminal;
	output [8:0] state;
	
	reg [8:0] state;
	reg odd, even, terminal;
	
	parameter  FIRST = 	9'b011_010_010;
	parameter  SECOND = 	9'b101_100_001;
	parameter  THIRD =	 	9'b010_111_010;
	parameter  FOURTH = 	9'b110_011_001;
	parameter  FIFTH = 	9'b101_010_110;
	
	always @(posedge clk or posedge rst) begin
		if (rst) state <= FIRST;
		else begin
			case (state)
				FIRST: 
					if (restart|pause) state <= FIRST;
					else state <= SECOND;
				SECOND: 
					if (restart) state <= FIRST;
					else if (pause) state <= SECOND;
					else state <= THIRD;
				THIRD:
					if (restart) state <= FIRST;
					else if (pause) state <= THIRD;
					else state <= FOURTH ;
				FOURTH:
					if (restart) state <= FIRST;
					else if (pause) state <= FOURTH;
					else state <= FIFTH;
				FIFTH:
					if (goto_third) state <= THIRD;
					else if (restart) state <= FIRST;
					else state <= FIFTH;
				
				default: state <= FIRST;
			endcase
		end
	end
	
	always @(*) begin
		odd = state[1];
		even = state[0];
		terminal = state[2];
		Out1 = state[8:6];
		Out2 = state[5:3];
	end
	
endmodule
				
					
	
